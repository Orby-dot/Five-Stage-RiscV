module pd
#(parameter  MEM_DEPTH = 32'd1048576)
(
  input clock,
  input reset
);

endmodule
